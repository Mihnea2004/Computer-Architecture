library verilog;
use verilog.vl_types.all;
entity counter_tb is
end counter_tb;
