library verilog;
use verilog.vl_types.all;
entity text2nibble_tb is
end text2nibble_tb;
