library verilog;
use verilog.vl_types.all;
entity cmp2b_tb is
end cmp2b_tb;
