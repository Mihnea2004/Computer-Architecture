library verilog;
use verilog.vl_types.all;
entity mul5bcd_tb is
end mul5bcd_tb;
