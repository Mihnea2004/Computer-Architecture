library verilog;
use verilog.vl_types.all;
entity seq3b_tb is
end seq3b_tb;
