library verilog;
use verilog.vl_types.all;
entity pktmux_tb is
end pktmux_tb;
