library verilog;
use verilog.vl_types.all;
entity msd_tb is
end msd_tb;
